/* Albert Wang (albertwa) & Tahmid Ahamed (ahamedt) */

`timescale 1ns / 1ps

// disable implicit wire declaration
`default_nettype none

module lc4_processor
   (input  wire        clk,                // main clock
    input wire         rst, // global reset
    input wire         gwe, // global we for single-step clock
                                    
    output wire [15:0] o_cur_pc, // Address to read from instruction memory
    input wire [15:0]  i_cur_insn, // Output of instruction memory
    output wire [15:0] o_dmem_addr, // Address to read/write from/to data memory
    input wire [15:0]  i_cur_dmem_data, // Output of data memory
    output wire        o_dmem_we, // Data memory write enable
    output wire [15:0] o_dmem_towrite, // Value to write to data memory
   
    output wire [1:0]  test_stall, // Testbench: is this is stall cycle? (don't compare the test values)
    output wire [15:0] test_cur_pc, // Testbench: program counter
    output wire [15:0] test_cur_insn, // Testbench: instruction bits
    output wire        test_regfile_we, // Testbench: register file write enable
    output wire [2:0]  test_regfile_wsel, // Testbench: which register to write in the register file 
    output wire [15:0] test_regfile_data, // Testbench: value to write into the register file
    output wire        test_nzp_we, // Testbench: NZP condition codes write enable
    output wire [2:0]  test_nzp_new_bits, // Testbench: value to write to NZP bits
    output wire        test_dmem_we, // Testbench: data memory write enable
    output wire [15:0] test_dmem_addr, // Testbench: address to read/write memory
    output wire [15:0] test_dmem_data, // Testbench: value read/writen from/to memory

    input wire [7:0]   switch_data, // Current settings of the Zedboard switches
    output wire [7:0]  led_data // Which Zedboard LEDs should be turned on?
    );

   
   
   /*** YOUR CODE HERE ***/

   /* Add $display(...) calls in the always block below to
    * print out debug information at the end of every cycle.
    * 
    * You may also use if statements inside the always block
    * to conditionally print out information.
    *
    * You do not need to resynthesize and re-implement if this is all you change;
    * just restart the simulation.
    */


    //F Stage
    assign led_data = switch_data;
    wire [15:0]   PC;
    wire [15:0]   next_pc;
    wire [15:0]   pcplusOne;

    cla16 add_one_to_pc(.a(PC), .b(16'b1), .cin(1'b0), .sum(pcplusOne));
    Nbit_reg #(16, 16'h8200) pc_reg_fetch_stage (.in(next_pc), .out(PC), .clk(clk), .we(1'b1), .gwe(gwe), .rst(rst));



    //D Stage
    wire [15:0]   decode_PC;
    Nbit_reg #(16, 16'h8200) pc_reg_decode_stage (.in(PC), .out(decode_PC), .clk(clk), .we(1'b1), .gwe(gwe), .rst(rst));

    wire [15:0]   decode_stage_instruction_output;
    Nbit_reg #(16, 16'd0) instruction_reg_decode_stage (.in(i_cur_insn), .out(decode_stage_instruction_output), .clk(clk), .we(1'b1), .gwe(gwe), .rst(rst));

    wire r1re;
    wire r2re;
    wire regfile_we;
    wire nzp_we;
    wire plus_one_select;
    wire is_load;
    wire is_store;
    wire is_branch;
    wire is_control_insn;

    wire [2:0]    r1_select;
    wire [2:0]    r2_select;
    wire [2:0]    rd_select;

    wire [15:0]   rsData;
    wire [15:0]   rtData;
    wire [15:0]   writeRegData;

    lc4_regfile decoder_regfile (
      .clk(clk),
      .gwe(gwe),
      .rst(rst),
      .i_rs(r1_select),
      .o_rs_data(rsData)
      .i_rt(r2_select),
      .o_rt_data(rtData),
      .i_rd(rd_select),
      .i_wdata(writeRegData),
      .i_rd_we(regfile_we)
    );

    lc4_decoder #(16) decoder(.insn(decode_stage_instruction_output), 
    .r1sel(r1_select), 
    .r1re(r1re), 
    .r2sel(r2_select),
    .wsel(rd_select),
    .regfile_we(regfile_we),
    .nzp_we(nzp_we),
    .select_pc_plus_one(plus_one_select),
    .is_load(is_load),
    .is_store(is_store),
    .is_branch(is_branch),
    .is_control_insn(is_control_insn)
    );
    
   
    //X Stage
    wire [15:0] x_PC;
    wire [15:0] x_stage_instruction_output;
    Nbit_reg #(16, 16'h8200) pc_reg_x_stage(.in(decode_PC), .out(x_PC), .clk(clk), .we(1'b1), .gwe(gwe), .rst(rst));
    Nbit_reg #(16, 16'd0) instruction_reg_execute_stage(.in(decode_stage_instruction_output), .out(x_stage_instruction_output), .clk(clk), .we(1'b1), .gwe(gwe), .rst(rst));
    Nbit_reg #(16, 16'd0) x_stage_write_data_reg
    Nbit_reg #(16, 16'd0) x_stage_rt_data_reg;
    Nbit_reg #(16, 16'd0) x_stage_rs_data_reg;


    //M Stage

    //W Stage



    //Test Wires
    assign o_cur_pc = PC;

`ifndef NDEBUG
   always @(posedge gwe) begin
      // $display("%d %h %h %h %h %h", $time, f_pc, d_pc, e_pc, m_pc, test_cur_pc);
      // if (o_dmem_we)
      //   $display("%d STORE %h <= %h", $time, o_dmem_addr, o_dmem_towrite);

      // Start each $display() format string with a %d argument for time
      // it will make the output easier to read.  Use %b, %h, and %d
      // for binary, hex, and decimal output of additional variables.
      // You do not need to add a \n at the end of your format string.
      // $display("%d ...", $time);

      // Try adding a $display() call that prints out the PCs of
      // each pipeline stage in hex.  Then you can easily look up the
      // instructions in the .asm files in test_data.

      // basic if syntax:
      // if (cond) begin
      //    ...;
      //    ...;
      // end

      // Set a breakpoint on the empty $display() below
      // to step through your pipeline cycle-by-cycle.
      // You'll need to rewind the simulation to start
      // stepping from the beginning.

      // You can also simulate for XXX ns, then set the
      // breakpoint to start stepping midway through the
      // testbench.  Use the $time printouts you added above (!)
      // to figure out when your problem instruction first
      // enters the fetch stage.  Rewind your simulation,
      // run it for that many nano-seconds, then set
      // the breakpoint.

      // In the objects view, you can change the values to
      // hexadecimal by selecting all signals (Ctrl-A),
      // then right-click, and select Radix->Hexadecimal.

      // To see the values of wires within a module, select
      // the module in the hierarchy in the "Scopes" pane.
      // The Objects pane will update to display the wires
      // in that module.

      //$display(); 
   end
`endif
endmodule
